module main

import txtar

fn main() {
}
